module inst_mem(
  output [31:0]	imem_instruction,
  input  clk,
  input  [31:0] imem_pc
);
  reg [31:0] cmd [256:0];
  reg [31:0] new_instruction;
  assign imem_instruction = new_instruction;
  initial begin
	// addi $t0, $0, 10
	cmd[4] <= 32'b00100000000010000000000000001010;
	// addi $t1, $0, 5
	cmd[8] <= 32'b00100000000010010000000000000101;
	// add $t2, $t1, $t0
	cmd[12] <= 32'b00000001001010000101000000100000;
	// add $t1, $t2, $t0
	cmd[16] <= 32'b00000001010010000100100000100000;
	// addi $t1, $t1, 20
	cmd[20] <= 32'b00100001001010010000000000010100;
	// add $t0, $t1, $t2
	cmd[24] <= 32'b00000001001010100100000000100000;
	// add $t1, $t0, $t2
	cmd[28] <= 32'b00000001000010100100100000100000;
	// add $t2, $t0, $t1
	cmd[32] <= 32'b00000001000010010101000000100000;
	// addi $t0, $t2, 10
	cmd[36] <= 32'b00100001010010000000000000001010;
	// addi $t2, $t2, 10
	cmd[40] <= 32'b00100001010010100000000000001010;
	// add $t2, $t2, $t0
	cmd[44] <= 32'b00000001010010000101000000100000;
	// slt $t3, $t0, $t2
	cmd[48] <= 32'b00000001000010100101100000101010;
	// slt $t3, $t2, $t0
	cmd[52] <= 32'b00000001010010000101100000101010;
	// sub $t2, $t1, $t0
	cmd[56] <= 32'b00000001001010000101000000100010;
	// addi $t2, $t2, 80
	cmd[60] <= 32'b00100001010010100000000001010000;
	// or $t3, $t0, $t1
	cmd[64] <= 32'b00000001000010010101100000100101;
	// and $t3, $t0, $t1
	cmd[68] <= 32'b00000001000010010101100000100100;
	// slti $t3, $t2, 15
	cmd[72] <= 32'b00101001010010110000000000001111;
	// addi $t0, $0, 10
	cmd[76] <= 32'b00100000000010000000000000001010;
	// sw $t0, 0($t0)
	cmd[80] <= 32'b10101101000010000000000000000000;
	// lw $t1, 0($t0)
	cmd[84] <= 32'b10001101000010010000000000000000;
  	// addi $t0, $0, 6
	cmd[88] <= 32'b00100000000010000000000000000110;
	// lw $t1, 4($t0)
	cmd[92] <= 32'b10001101000010010000000000000100;
	// sw $t1, 1($t0)
	cmd[96] <= 32'b10101101000010010000000000000001;
	// sw $t1, 2($t0)
	cmd[100] <= 32'b10101101000010010000000000000010;
	// lw $t0, 1($t0)
	cmd[104] <= 32'b10001101000010000000000000000001;
	// lw $t2, 2($t0)
	cmd[108] <= 32'b10001101000010100000000000000001;
	// addi $t0, $0, 15
	cmd[112] <= 32'b00100000000010000000000000001111;
	// addi $t1, $0, 15
	cmd[116] <= 32'b00100000000010010000000000001111;
	// beq $t0, $t1, 4
	cmd[120] <= 32'b00010001000010010000000000000100;
	// Test for beq
	cmd[124] <= 32'bx;
	cmd[128] <= 32'bx;
	cmd[132] <= 32'bx;
	cmd[136] <= 32'bx;
	// j -35 : reset to begin
	cmd[140] <= 32'b00001011111111111111111111011101;
  end
  always @(imem_pc) begin
	new_instruction[31:0] = cmd[imem_pc][31:0];
  end

endmodule 
